Library ieee;
Use ieee.std_logic_1164.all;

ENTITY ForwardingUnit IS

PORT(
	Reset: IN std_logic;
	
	ID_EX_RS1,ID_EX_RS2,ID_EX_RD: IN std_logic_vector (2 DOWNTO 0);
	ID_EX_SOURCECONTROL: IN std_logic_vector(2 DOWNTO 0);
	EX_MEM_RS1,EX_MEM_RD: IN std_logic_vector (2 DOWNTO 0);
	EX_MEM_DSTCONTROL: IN std_logic_vector (1 DOWNTO 0);
	MEM_WB_RS1,MEM_WB_RD: IN std_logic_vector (2 DOWNTO 0);
	MEM_WB_DSTCONTROL: IN std_logic_vector (1 DOWNTO 0);
	REG_WRITE_EX_MEM: IN std_logic;
	REG_WRITE_MEM_WB: IN std_logic;
	RS1_SELECT: OUT std_logic_vector (2 downto 0);
	RS2_SELECT: OUT std_logic_vector (2 downto 0);
	RD_SELECT: OUT std_logic_vector (2 downto 0)
	
);
	
end ForwardingUnit;

ARCHITECTURE a_ForwardingUnit of ForwardingUnit 
IS
	SIGNAL RS1_SELECT_MEM,RS2_SELECT_MEM,RD_SELECT_MEM: std_logic;
	SIGNAL RS1_SELECT_WB,RS2_SELECT_WB,RD_SELECT_WB: std_logic;
Begin


	RS1_SELECT_MEM <= '1' WHEN (ID_EX_SOURCECONTROL = "001") and (EX_MEM_DSTCONTROL = "01") and (ID_EX_RS1 = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "001") and (EX_MEM_DSTCONTROL = "10") and (ID_EX_RS1 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "001") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS1 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "001") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS1 = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "01") and (ID_EX_RS1 = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "10") and (ID_EX_RS1 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS1 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS1 = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "01") and (ID_EX_RS1 = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "10") and (ID_EX_RS1 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS1 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS1 = EX_MEM_RD)
	ELSE '0';

	RS1_SELECT_WB <= '1' WHEN (ID_EX_SOURCECONTROL = "001") and (MEM_WB_DSTCONTROL = "01") and (ID_EX_RS1 = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "001") and (MEM_WB_DSTCONTROL = "10") and (ID_EX_RS1 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "001") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS1 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "001") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS1 = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "01") and (ID_EX_RS1 = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "10") and (ID_EX_RS1 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS1 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS1 = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "01") and (ID_EX_RS1 = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "10") and (ID_EX_RS1 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS1 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS1 = MEM_WB_RD)
	ELSE '0';




	RS2_SELECT_MEM <= '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "01") and (ID_EX_RS2 = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "10") and (ID_EX_RS2 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS2 = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RS2 = EX_MEM_RD)
	ELSE '0';

	RS2_SELECT_WB <= '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "01") and (ID_EX_RS2 = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "10") and (ID_EX_RS2 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS2 = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "100") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RS2 = MEM_WB_RD)
	ELSE '0';


	RD_SELECT_MEM <= '1' WHEN (ID_EX_SOURCECONTROL = "010") and (EX_MEM_DSTCONTROL = "01") and (ID_EX_RD = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "010") and (EX_MEM_DSTCONTROL = "10") and (ID_EX_RD = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "010") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RD = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "010") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RD = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "01") and (ID_EX_RD = EX_MEM_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "10") and (ID_EX_RD = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RD = EX_MEM_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (EX_MEM_DSTCONTROL = "11") and (ID_EX_RD = EX_MEM_RD)
	ELSE '0';

	RD_SELECT_WB <= '1' WHEN (ID_EX_SOURCECONTROL = "010") and (MEM_WB_DSTCONTROL = "01") and (ID_EX_RD = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "010") and (MEM_WB_DSTCONTROL = "10") and (ID_EX_RD = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "010") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RD = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "010") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RD = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "01") and (ID_EX_RD = MEM_WB_RD)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "10") and (ID_EX_RD = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RD = MEM_WB_RS1)
	ELSE '1' WHEN (ID_EX_SOURCECONTROL = "111") and (MEM_WB_DSTCONTROL = "11") and (ID_EX_RD = MEM_WB_RD)
	ELSE '0';


	RS1_SELECT <= "001" WHEN RS1_SELECT_MEM = '0' AND RS1_SELECT_WB = '0'
	ELSE "010" WHEN RS1_SELECT_MEM = '1'
	ELSE "100" WHEN RS1_SELECT_WB = '1';
	
	RS2_SELECT <= "001" WHEN RS2_SELECT_MEM ='0' AND RS2_SELECT_WB ='0'
	ELSE "010" WHEN RS2_SELECT_MEM = '1'
	ELSE "100" WHEN RS2_SELECT_WB = '1';

	RD_SELECT <= "001" WHEN RD_SELECT_MEM = '0' AND RD_SELECT_WB = '0'
	ELSE "010" WHEN RD_SELECT_MEM ='1'
	ELSE "100" WHEN RD_SELECT_WB = '1';




END a_ForwardingUnit;


